module VGA_pic(
input wire vga_clk , //输入工作时钟,频率25MHz
input wire sys_rst_n , //输入复位信号,低电平有效
input wire [9:0] pix_x , //输入有效显示区域像素点X轴坐标
input wire [9:0] pix_y , //输入有效显示区域像素点Y轴坐标

output reg [15:0] pix_data //输出像素点色彩信息

);

////
//\* Parameter and Internal Signal \//
////
//parameter define
parameter CHAR_B_H= 10'd192 , //字符开始X轴坐标
CHAR_B_V= 10'd208 ; //字符开始Y轴坐标

parameter CHAR_W = 10'd256 , //字符宽度
CHAR_H = 10'd64 ; //字符高度

parameter BLACK = 16'h0000, //黑色
WHITE = 16'hFFFF, //白色
GOLDEN = 16'hFEC0; //金色

//wire define
wire [9:0] char_x ; //字符显示X轴坐标
wire [9:0] char_y ; //字符显示Y轴坐标

//reg define
reg [255:0] char [63:0] ; //字符数据

////
//\* Main Code \//
////

//字符显示坐标
assign char_x = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
? (pix_x - CHAR_B_H) : 10'h3FF;
assign char_y = (((pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W)))
&&((pix_y >= CHAR_B_V)&&(pix_y < (CHAR_B_V + CHAR_H))))
? (pix_y - CHAR_B_V) : 10'h3FF;

//char:字符数据
always@(posedge vga_clk)
begin
 char [0] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
 char [1] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
 char [2] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
 char [3] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
 char [4] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
 char [5] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
 char [6] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
 char [7] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
 char [8] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
 char [9] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
char [10] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
char [11] <= 63'h0000FF8003FF000000007FF807FE00000000001FE000000000000FFFFFF00000;
char [12] <= 63'h0000FF8003FF000000007FF807FE00000000007FF880000000000FFFFFF00000;
char [13] <= 63'h00001F8003F8000000000FC000F00000000000F03F80000000000F03C0F80000;
char [14] <= 63'h00001F8003F800000000078000600000000001C00F80000000001E03C0380000;
char [15] <= 63'h00001F8007F800000000078000600000000003C00780000000001C03C0380000;
char [16] <= 63'h00001FC007F8000000000780006000000000078003C0000000001803C0180000;
char [17] <= 63'h00001FC007F8000000000780006000000000078001C0000000001803C0180000;
char [18] <= 63'h00001FC007F8000000000780006000000000070001C0000000001003C00C0000;
char [19] <= 63'h00001FC00FF80000000007800060000000000F0000C0000000003003C00C0000;
char [20] <= 63'h00001FE00FF80000000007800060000000000F0000C0000000003003C0040000;
char [21] <= 63'h00001FE00FF80000000007800060000000000F000000000000000003C0000000;
char [22] <= 63'h00001FE00FF80000000007800060000000000F000000000000000003C0000000;
char [23] <= 63'h00001FE00FF80000000007800060000000000F000000000000000003C0000000;
char [24] <= 63'h00001FE01FF80000000007800060000000000F800000000000000003C0000000;
char [25] <= 63'h00001FF01FF800000000078000600000000007C00000000000000003C0000000;
char [26] <= 63'h00001FF01DF800000000078000600000000007E00000000000000003C0000000;
char [27] <= 63'h00001DF01DF800000000078000600000000007F00000000000000003C0000000;
char [28] <= 63'h00001DF03DF800000000078000600000000003FC0000000000000003C0000000;
char [29] <= 63'h00001DF83DF800000000078000600000000001FF0000000000000003C0000000;
char [30] <= 63'h00001DF839F8000000000780006000000000007FC000000000000003C0000000;
char [31] <= 63'h00001CF839F8000000000780006000000000003FF000000000000003C0000000;
char [32] <= 63'h00001CF879F8000000000780006000000000000FFC00000000000003C0000000;
char [33] <= 63'h00001CF879F80000000007800060000000000003FE00000000000003C0000000;
char [34] <= 63'h00001CFC71F80000000007800060000000000000FF00000000000003C0000000;
char [35] <= 63'h00001C7C71F800000000078000600000000000003F80000000000003C0000000;
char [36] <= 63'h00001C7CF1F800000000078000600000000000000FC0000000000003C0000000;
char [37] <= 63'h00001C7CF1F8000000000780006000000000000007E0000000000003C0000000;
char [38] <= 63'h00001C7EE1F8000000000780006000000000000003E0000000000003C0000000;
char [39] <= 63'h00001C7EE1F8000000000780006000000000000001E0000000000003C0000000;
char [40] <= 63'h00001C3EE1F8000000000780006000000000000001F0000000000003C0000000;
char [41] <= 63'h00001C3FE1F8000000000780006000000000000000F0000000000003C0000000;
char [42] <= 63'h00001C3FE1F8000000000780006000000000080000F0000000000003C0000000;
char [43] <= 63'h00001C3FC1F8000000000780006000000000180000F0000000000003C0000000;
char [44] <= 63'h00001C1FC1F8000000000780006000000000180000F0000000000003C0000000;
char [45] <= 63'h00001C1FC1F80000000007800060000000001C0000F0000000000003C0000000;
char [46] <= 63'h00001C1FC1F80000000007800060000000000C0000F0000000000003C0000000;
char [47] <= 63'h00001C1F81F800000000078000E0000000000E0000E0000000000003C0000000;
char [48] <= 63'h00001C1F81F800000000038000C0000000000E0001E0000000000003C0000000;
char [49] <= 63'h00001C0F81F80000000003C001C0000000000F0001C0000000000003C0000000;
char [50] <= 63'h00001C0F81F80000000001C00380000000000F8003C0000000000003C0000000;
char [51] <= 63'h00001C0F01F80000000001E00700000000000FC00780000000000003C0000000;
char [52] <= 63'h0000FF8F0FFF0000000000F81E000000000007F81F00000000000007E0000000;
char [53] <= 63'h0000FF870FFF00000000003FFC0000000000061FFC0000000000007FFE000000;
char [54] <= 63'h00000000000000000000000FE000000000000407F00000000000007FFE000000;
char [55] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
char [56] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
char [57] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
char [58] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
char [59] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
char [60] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
char [61] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
char [62] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
char [63] <= 63'h0000000000000000000000000000000000000000000000000000000000000000;
 end

 //pix_data:输出像素点色彩信息,根据当前像素点坐标指定当前像素点颜色数据
 always@(posedge vga_clk or negedge sys_rst_n)
 if(sys_rst_n == 1'b0)
 pix_data <= BLACK;
 else if((((pix_x >= (CHAR_B_H - 1'b1))
 && (pix_x < (CHAR_B_H + CHAR_W -1'b1)))
 && ((pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H))))
 && (char[char_y][10'd255 - char_x] == 1'b1))
 pix_data <= GOLDEN;
 else
 pix_data <= BLACK;

 endmodule